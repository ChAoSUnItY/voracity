module main

import voracity.complete.bytes
import voracity.complete.character

fn main() {
}

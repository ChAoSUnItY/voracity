module main

import voracity.complete.bytes
import voracity.complete.character

fn main() {
	println(typeof[character.CharParser]())
	println(typeof[character.CharParserOpt]())
}

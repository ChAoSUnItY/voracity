module main

import voracity

fn main() {
	println('Hello World!')
}

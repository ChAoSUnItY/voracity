module tests

fn test_alt() {

}

module voracity

type VoidParser = fn (mut State)
